version https://git-lfs.github.com/spec/v1
oid sha256:7a6ea0f48e48fbf400afb0ab51b0f0b370b914c3f06b4c70fd9eb99a71238b21
size 104858112
